module bin16_to_bcd(output reg [3:0] digit [0:4], input [15:0] bin);
    
endmodule
