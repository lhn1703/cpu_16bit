module test1(output a);
	assign a = 1;
endmodule
