module cpu_16bit (output [15:0] result_reg, input [15:0] initial_input, input clk, pc_reset);
    
	// IF
	
	
	// IF/ID
	
	
	// ID
	
	
	// ID/EX
	
	
	// EX
	
	
	// EX/MEM
	
	
	// MEM
	
	
	// MEM/WB
	
	
	// WB
	
	
	// Pipelining

endmodule